��  CCircuit��  CSerializeHack           ��  CPart    H   H     ��� 	 CResistor��  CValue  � � $    10M       �cA      �?M  �� 	 CTerminal  � (� )               �          �  � (� )                            � $� ,        ��      ��  CEarth�  p 0q E                             c D{ L         ��      �� 	 CVoltRail
�  � � � �     3.2V(    ������	@      �? V �  � � � 	     
   ������	@wb:����    � � � �         ����     ��  CSPDT��  CToggle  � 8X        �  � T� i        ������	@wb:����  �  � (� =      
   ������	@wb:���>  �  � (� =                �            � <� T         ��    ��  �(�=                             �<�D         ��      �
�  h�    10M       �cA      �?M  �  � �!                          �  X m!     	          �            l�$    !    ��      �
�  � ;�     3.2V(    ������	@      �? V �  @� A�         ������	@�˦A���    <� D�     %    ����     �� 
 CPushBreak��  CKey  L� p      '   �  @A        ������	@�˦A���  �  @� A�        	 ������	@�˦A��>    <� F    *      ��    ��  X8xX      ,   �  HTIi        ������	@�˦A���  �  P(Q=      	          �          �  @(A=         ������	@�˦A��>    <<TT    .      ��    ��  � (� =                 tԖ��?    � <� D     2    ��      �� 
 CVoltmeter��  CMeter  �,�     3.18   �  $9	        ��_ido	@          �  � 	                            �$    7    ��      �
�  �(�    100k        j�@      �?k  �  $�9�        ��_ido	@o�˦A��>  �  � ��        �G�%;��?o�˦A���    �$�    ;    ��      �
�  � �� �    27k          ^�@      �?k  �  � �� �         �G�%;��?tԖ��?  �  � �� 	                tԖ���    � �� �     ?    ��      �
�  #�C�    1k          @�@      �?k  �  HhI}       	 ������	@�˦A��>  �  H�I�        ��_ido	@�˦A���    D|L�     C    ��      �
�  � �� �    100k          j�@      �?k  �  � h� }       	 ������	@wb:���>  �  � �� �        �G�%;��?wb:����    � |� �     G    ��          H   H     ���  CWire  H�I	       J�  H�I�       J�  � �� �       J�  � (� )      J�  p (q 1       J�  p (� )      J�  � � )      
 J�  � �)       J�  � �!      J�  P Q)      	 J�  P Y!     	 J�  @A)       J�  � � )       J�  8�I�      J�  8I	      J�  � � 	      J�  � �� �      J�  � �� �          H   H     �    H   H         H   H       N  P   O    Q   G  Q   N   R  ! ! S " U " % % + * * V + % + . . C / T / 0 V 0 2 W 2 7 7 Y 8 Z 8 ; ; X < [ < ? \ ? @ @ W C . C D D L G  G H H M X Y D K H [   P  O    S  ! R U / T " * 0 Z 2 ; L 7 K @ 8 \ < ? M            �$s�        @     +        @            @    "V  (      �h                
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 